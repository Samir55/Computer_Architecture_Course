library ieee;
use ieee.std_logic_1164.all;

-- MAR register module connected with read/write enable ready to be integrated in the control cicuit.
Entity MARRegister is 
	Generic (n: integer := 16);
	port(InternalBus: inout std_logic_vector(n-1 downTo 0); RamAddress: out std_logic_vector(n-1 downTo 0); Clk, Rst, WriteEnable, ReadEnable: in std_logic);
End Entity MARRegister;

Architecture MARRegisterImplementation of MARRegister is 

	Component nBitRegister is 
		Generic (n: integer := 16);
		port(D: in std_logic_vector(n-1 downTo 0); Q: out std_logic_vector(n-1 downTo 0); Clk, Rst: in std_logic);
	End Component;

	Component TriStateBuff is 
		Generic (n: integer := 16);
		port(A: in std_logic_vector(n-1 downTo 0); Enable: in std_logic; B: out std_logic_vector(n-1 downTo 0));
	End Component;
	
	Signal RegisterInputD, RegisterOutputQ: std_logic_vector(n-1 downTo 0);
Begin
	WriteTriStateBuffer: TriStateBuff GENERIC MAP (n=>16) PORT MAP(InternalBus, WriteEnable, RegisterInputD); -- Write Enable means write a value to this register.
	ReadTriStateBuffer: TriStateBuff GENERIC MAP (n=>16) PORT MAP(RegisterOutputQ, ReadEnable, InternalBus);
	NRegister : nBitRegister GENERIC MAP (n=>16) PORT MAP(RegisterInputD, RegisterOutputQ, Clk, Rst);
	RamAddress <= RegisterOutputQ;

End MARRegisterImplementation;




